module LDA_control (
	input clk,
	input reset,

	input i_start,
	
	// Datapath
	input i_done,
	output logic o_setup,
	output logic o_step
);



endmodule
