module LDA (
	input clk,
	input reset,

	input i_start,
	input [8:0] i_x0,
	input [7:0] i_y0,
	input [8:0] i_x1,
	input [7:0] i_y1,
	input [2:0] i_col,
	
	output o_done
);



endmodule
