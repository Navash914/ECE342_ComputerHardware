module LDA_datapath (
	input clk,
	input reset,
	
	input [8:0] i_x0,
	input [7:0] i_y0,
	input [8:0] i_x1,
	input [7:0] i_y1,
	
	input i_setup,
	input i_step
	
	output o_plot,
	output o_done
);



endmodule
