module UI_control (
	input clk,
	input reset,
	
	input i_go,
	input i_done,
	
	output o_start
);



endmodule
