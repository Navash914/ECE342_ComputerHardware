module asc_datapath (
	input clk,
	input reset,
	
	input [31:0] i_address,
	input [31:0] i_writedata,
	output [31:0] o_read_data
);



endmodule
